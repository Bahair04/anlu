module four_channel_video_splicer
#(
    parameter  integer                   AXI_DATA_WIDTH = 32,	//SDRAM����λ��
	parameter  integer                   AXI_ADDR_WIDTH = 21	//SDRAM��ַλ��
)(

);

endmodule